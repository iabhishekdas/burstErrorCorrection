module encoder (
	input [0:15] m,
	output [0:24] c
);

	wire [0:8] p;

	assign p[0] = m[0] ^ m[4] ^ m[8] ^ m[12];
	assign p[1] = m[1] ^ m[5] ^ m[9] ^ m[13];
	assign p[2] = m[2] ^ m[6] ^ m[10] ^ m[14];
	assign p[3] = m[3] ^ m[7] ^ m[11] ^ m[15];
	assign p[4] = m[0] ^ m[2] ^ m[6] ^ m[7] ^ m[8] ^ m[11];
	assign p[5] = m[0] ^ m[3] ^ m[6] ^ m[9] ^ m[12];
	assign p[6] = m[0] ^ m[1] ^ m[4] ^ m[6] ^ m[7] ^ m[10] ^ m[13];
	assign p[7] = m[0] ^ m[2] ^ m[3] ^ m[6] ^ m[7] ^ m[8] ^ m[9] ^ m[10] ^ m[14];
	assign p[8] = m[1] ^ m[2] ^ m[5] ^ m[6] ^ m[8] ^ m[9] ^ m[10] ^ m[11] ^ m[15];

	assign c = {m,p};

endmodule

module decoder (
	input [0:24] c,
	output [0:15] m
);

	wire [0:8] p, s;
	wire [0:15] b, en;
	assign b = c[0:15];
	assign p = c[16:24];

	assign s[0] = p[0] ^ b[0] ^ b[4] ^ b[8] ^ b[12];
	assign s[1] = p[1] ^ b[1] ^ b[5] ^ b[9] ^ b[13];
	assign s[2] = p[2] ^ b[2] ^ b[6] ^ b[10] ^ b[14];
	assign s[3] = p[3] ^ b[3] ^ b[7] ^ b[11] ^ b[15];
	assign s[4] = p[4] ^ b[0] ^ b[2] ^ b[6] ^ b[7] ^ b[8] ^ b[11];
	assign s[5] = p[5] ^ b[0] ^ b[3] ^ b[6] ^ b[9] ^ b[12];
	assign s[6] = p[6] ^ b[0] ^ b[1] ^ b[4] ^ b[6] ^ b[7] ^ b[10] ^ b[13];
	assign s[7] = p[7] ^ b[0] ^ b[2] ^ b[3] ^ b[6] ^ b[7] ^ b[8] ^ b[9] ^ b[10] ^ b[14];
	assign s[8] = p[8] ^ b[1] ^ b[2] ^ b[5] ^ b[6] ^ b[8] ^ b[9] ^ b[10] ^ b[11] ^ b[15];

	assign en[0] = (s[4] ^ s[0] ^ s[2]) | (s[5] ^ s[0] ^ s[3]) | (s[6] ^ s[0] ^ s[1]) | (s[7] ^ s[0] ^ s[2] ^ s[3]) | (s[8] ^ s[1] ^ s[2]);
	assign en[1] = (s[4] ^ s[2]) | (s[5] ^ s[3]) | (s[6] ^ s[1] ^ s[0]) | (s[7] ^ s[2] ^ s[3]) | (s[8] ^ s[1] ^ s[2]);
	assign en[2] = (s[4] ^ s[2]) | (s[5] ^ s[3]) | (s[6] ^ s[0]) | (s[7] ^ s[2] ^ s[3]) | (s[8] ^ s[2] ^ s[1]);
	assign en[3] = (s[4] ^ s[2]) | (s[5] ^ s[3] ^ s[2]) | (s[6] ^ s[0] ^ s[2]) | (s[7] ^ s[3] ^ s[2]) | (s[8] ^ s[1] ^ s[2]);
	assign en[4] = (s[4] ^ s[2] ^ s[3]) | (s[5] ^ s[2]) | (s[6] ^ s[0] ^ s[2] ^ s[3]) | (s[7] ^ s[2] ^ s[3]) | (s[8] ^ s[1] ^ s[2]);
	assign en[5] = (s[4] ^ s[2] ^ s[3] ^ s[0]) | (s[5] ^ s[2]) | (s[6] ^ s[2] ^ s[3]) | (s[7] ^ s[2] ^ s[3] ^ s[0]) | (s[8] ^ s[1] ^ s[2] ^ s[0]);
	assign en[6] = (s[4] ^ s[2] ^ s[3] ^ s[0]) | (s[5] ^ s[2] ^ s[1]) | (s[6] ^ s[2] ^ s[3]) | (s[7] ^ s[2] ^ s[3] ^ s[0] ^ s[1]) | (s[8] ^ s[2] ^ s[0] ^ s[1]);
	assign en[7] = (s[4] ^ s[3] ^ s[0]) | (s[5] ^ s[1]) | (s[6] ^ s[3] ^ s[2]) | (s[7] ^ s[3] ^ s[0] ^ s[1] ^ s[2]) | (s[8] ^ s[0] ^ s[1] ^ s[2]);
	assign en[8] = (s[4] ^ s[0] ^ s[3]) | (s[5] ^ s[1]) | (s[6] ^ s[2]) | (s[7] ^ s[0] ^ s[1] ^ s[2]) | (s[8] ^ s[0] ^ s[1] ^ s[2] ^ s[3]);
	assign en[9] = (s[4] ^ s[3]) | (s[5] ^ s[1] ^ s[0]) | (s[6] ^ s[2]) | (s[7] ^ s[1] ^ s[2]) | (s[8] ^ s[1] ^ s[2] ^ s[3]);
	assign en[10] = (s[4] ^ s[3]) | (s[5] ^ s[0]) | (s[6] ^ s[2] ^ s[1]) | (s[7] ^ s[2]) | (s[8] ^ s[2] ^ s[3]);
	assign en[11] = (s[4] ^ s[3]) | (s[5] ^ s[0]) | (s[6] ^ s[1]) | (s[7] ^ s[2]) | (s[8] ^ s[3]);
	assign en[12] = (s[4]) | (s[5] ^ s[0]) | (s[6] ^ s[1]) | (s[7] ^ s[2]) | (s[8] ^ s[3]);
	assign en[13] = (s[4]) | (s[5]) | (s[6] ^ s[1]) | (s[7] ^ s[2]) | (s[8] ^ s[3]);
	assign en[14] = (s[4]) | (s[5]) | (s[6]) | (s[7] ^ s[2]) | (s[8] ^ s[3]);
	assign en[15] = (s[4]) | (s[5]) | (s[6]) | (s[7]) | (s[8] ^ s[3]);

	assign m[0] = ((~( en[0] )) & s[0]) ^ b[0];
	assign m[1] = ((~( en[1] & en[0] )) & s[1]) ^ b[1];
	assign m[2] = ((~( en[2] & en[1] & en[0] )) & s[2]) ^ b[2];
	assign m[3] = ((~( en[3] & en[2] & en[1] & en[0] )) & s[3]) ^ b[3];
	assign m[4] = ((~( en[4] & en[3] & en[2] & en[1] )) & s[0]) ^ b[4];
	assign m[5] = ((~( en[5] & en[4] & en[3] & en[2] )) & s[1]) ^ b[5];
	assign m[6] = ((~( en[6] & en[5] & en[4] & en[3] )) & s[2]) ^ b[6];
	assign m[7] = ((~( en[7] & en[6] & en[5] & en[4] )) & s[3]) ^ b[7];
	assign m[8] = ((~( en[8] & en[7] & en[6] & en[5] )) & s[0]) ^ b[8];
	assign m[9] = ((~( en[9] & en[8] & en[7] & en[6] )) & s[1]) ^ b[9];
	assign m[10] = ((~( en[10] & en[9] & en[8] & en[7] )) & s[2]) ^ b[10];
	assign m[11] = ((~( en[11] & en[10] & en[9] & en[8] )) & s[3]) ^ b[11];
	assign m[12] = ((~( en[12] & en[11] & en[10] & en[9] )) & s[0]) ^ b[12];
	assign m[13] = ((~( en[13] & en[12] & en[11] & en[10] )) & s[1]) ^ b[13];
	assign m[14] = ((~( en[14] & en[13] & en[12] & en[11] )) & s[2]) ^ b[14];
	assign m[15] = ((~( en[15] & en[14] & en[13] & en[12] )) & s[3]) ^ b[15];

endmodule