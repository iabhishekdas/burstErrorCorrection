module encoder (
	input [0:63] m,
	output [0:74] c
);

	wire [0:10] p;

	assign p[0] = m[0] ^ m[4] ^ m[8] ^ m[12] ^ m[16] ^ m[20] ^ m[24] ^ m[28] ^ m[32] ^ m[36] ^ m[40] ^ m[44] ^ m[48] ^ m[52] ^ m[56] ^ m[60];
	assign p[1] = m[1] ^ m[5] ^ m[9] ^ m[13] ^ m[17] ^ m[21] ^ m[25] ^ m[29] ^ m[33] ^ m[37] ^ m[41] ^ m[45] ^ m[49] ^ m[53] ^ m[57] ^ m[61];
	assign p[2] = m[2] ^ m[6] ^ m[10] ^ m[14] ^ m[18] ^ m[22] ^ m[26] ^ m[30] ^ m[34] ^ m[38] ^ m[42] ^ m[46] ^ m[50] ^ m[54] ^ m[58] ^ m[62];
	assign p[3] = m[3] ^ m[7] ^ m[11] ^ m[15] ^ m[19] ^ m[23] ^ m[27] ^ m[31] ^ m[35] ^ m[39] ^ m[43] ^ m[47] ^ m[51] ^ m[55] ^ m[59] ^ m[63];
	assign p[4] = m[1] ^ m[4] ^ m[8] ^ m[15] ^ m[16] ^ m[18] ^ m[19] ^ m[22] ^ m[25] ^ m[28] ^ m[29] ^ m[30] ^ m[31] ^ m[33] ^ m[34] ^ m[35] ^ m[40] ^ m[41] ^ m[42] ^ m[43] ^ m[52] ^ m[53] ^ m[54] ^ m[55];
	assign p[5] = m[5] ^ m[6] ^ m[8] ^ m[10] ^ m[11] ^ m[14] ^ m[15] ^ m[16] ^ m[17] ^ m[20] ^ m[26] ^ m[28] ^ m[30] ^ m[32] ^ m[33] ^ m[34] ^ m[36] ^ m[37] ^ m[40] ^ m[44] ^ m[45] ^ m[46] ^ m[47] ^ m[52] ^ m[56] ^ m[57] ^ m[58];
	assign p[6] = m[1] ^ m[5] ^ m[7] ^ m[9] ^ m[10] ^ m[14] ^ m[15] ^ m[18] ^ m[21] ^ m[23] ^ m[28] ^ m[29] ^ m[30] ^ m[31] ^ m[32] ^ m[36] ^ m[38] ^ m[39] ^ m[41] ^ m[44] ^ m[48] ^ m[49] ^ m[53] ^ m[59];
	assign p[7] = m[0] ^ m[5] ^ m[6] ^ m[9] ^ m[12] ^ m[14] ^ m[15] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[20] ^ m[21] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[29] ^ m[30] ^ m[31] ^ m[32] ^ m[33] ^ m[36] ^ m[37] ^ m[38] ^ m[39] ^ m[41] ^ m[42] ^ m[45] ^ m[48] ^ m[50] ^ m[54] ^ m[60];
	assign p[8] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[7] ^ m[8] ^ m[9] ^ m[14] ^ m[15] ^ m[16] ^ m[17] ^ m[19] ^ m[20] ^ m[21] ^ m[28] ^ m[29] ^ m[31] ^ m[32] ^ m[34] ^ m[35] ^ m[36] ^ m[37] ^ m[38] ^ m[42] ^ m[44] ^ m[46] ^ m[48] ^ m[50] ^ m[51] ^ m[56] ^ m[61];
	assign p[9] = m[0] ^ m[2] ^ m[5] ^ m[6] ^ m[7] ^ m[11] ^ m[12] ^ m[14] ^ m[16] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[24] ^ m[27] ^ m[28] ^ m[29] ^ m[33] ^ m[35] ^ m[37] ^ m[38] ^ m[39] ^ m[40] ^ m[43] ^ m[47] ^ m[49] ^ m[50] ^ m[51] ^ m[55] ^ m[57] ^ m[62];
	assign p[10] = m[0] ^ m[1] ^ m[2] ^ m[3] ^ m[6] ^ m[7] ^ m[13] ^ m[14] ^ m[17] ^ m[18] ^ m[20] ^ m[22] ^ m[23] ^ m[24] ^ m[25] ^ m[27] ^ m[29] ^ m[30] ^ m[31] ^ m[32] ^ m[34] ^ m[35] ^ m[39] ^ m[43] ^ m[45] ^ m[46] ^ m[47] ^ m[49] ^ m[51] ^ m[58] ^ m[59] ^ m[63];

	assign c = {m,p};

endmodule

module decoder (
	input [0:74] c,
	output [0:63] m
);

	wire [0:10] p, s;
	wire [0:63] b, en;
	assign b = c[0:63];
	assign p = c[64:74];

	assign s[0] = p[0] ^ b[0] ^ b[4] ^ b[8] ^ b[12] ^ b[16] ^ b[20] ^ b[24] ^ b[28] ^ b[32] ^ b[36] ^ b[40] ^ b[44] ^ b[48] ^ b[52] ^ b[56] ^ b[60];
	assign s[1] = p[1] ^ b[1] ^ b[5] ^ b[9] ^ b[13] ^ b[17] ^ b[21] ^ b[25] ^ b[29] ^ b[33] ^ b[37] ^ b[41] ^ b[45] ^ b[49] ^ b[53] ^ b[57] ^ b[61];
	assign s[2] = p[2] ^ b[2] ^ b[6] ^ b[10] ^ b[14] ^ b[18] ^ b[22] ^ b[26] ^ b[30] ^ b[34] ^ b[38] ^ b[42] ^ b[46] ^ b[50] ^ b[54] ^ b[58] ^ b[62];
	assign s[3] = p[3] ^ b[3] ^ b[7] ^ b[11] ^ b[15] ^ b[19] ^ b[23] ^ b[27] ^ b[31] ^ b[35] ^ b[39] ^ b[43] ^ b[47] ^ b[51] ^ b[55] ^ b[59] ^ b[63];
	assign s[4] = p[4] ^ b[1] ^ b[4] ^ b[8] ^ b[15] ^ b[16] ^ b[18] ^ b[19] ^ b[22] ^ b[25] ^ b[28] ^ b[29] ^ b[30] ^ b[31] ^ b[33] ^ b[34] ^ b[35] ^ b[40] ^ b[41] ^ b[42] ^ b[43] ^ b[52] ^ b[53] ^ b[54] ^ b[55];
	assign s[5] = p[5] ^ b[5] ^ b[6] ^ b[8] ^ b[10] ^ b[11] ^ b[14] ^ b[15] ^ b[16] ^ b[17] ^ b[20] ^ b[26] ^ b[28] ^ b[30] ^ b[32] ^ b[33] ^ b[34] ^ b[36] ^ b[37] ^ b[40] ^ b[44] ^ b[45] ^ b[46] ^ b[47] ^ b[52] ^ b[56] ^ b[57] ^ b[58];
	assign s[6] = p[6] ^ b[1] ^ b[5] ^ b[7] ^ b[9] ^ b[10] ^ b[14] ^ b[15] ^ b[18] ^ b[21] ^ b[23] ^ b[28] ^ b[29] ^ b[30] ^ b[31] ^ b[32] ^ b[36] ^ b[38] ^ b[39] ^ b[41] ^ b[44] ^ b[48] ^ b[49] ^ b[53] ^ b[59];
	assign s[7] = p[7] ^ b[0] ^ b[5] ^ b[6] ^ b[9] ^ b[12] ^ b[14] ^ b[15] ^ b[16] ^ b[17] ^ b[18] ^ b[19] ^ b[20] ^ b[21] ^ b[22] ^ b[24] ^ b[26] ^ b[28] ^ b[29] ^ b[30] ^ b[31] ^ b[32] ^ b[33] ^ b[36] ^ b[37] ^ b[38] ^ b[39] ^ b[41] ^ b[42] ^ b[45] ^ b[48] ^ b[50] ^ b[54] ^ b[60];
	assign s[8] = p[8] ^ b[0] ^ b[2] ^ b[3] ^ b[5] ^ b[7] ^ b[8] ^ b[9] ^ b[14] ^ b[15] ^ b[16] ^ b[17] ^ b[19] ^ b[20] ^ b[21] ^ b[28] ^ b[29] ^ b[31] ^ b[32] ^ b[34] ^ b[35] ^ b[36] ^ b[37] ^ b[38] ^ b[42] ^ b[44] ^ b[46] ^ b[48] ^ b[50] ^ b[51] ^ b[56] ^ b[61];
	assign s[9] = p[9] ^ b[0] ^ b[2] ^ b[5] ^ b[6] ^ b[7] ^ b[11] ^ b[12] ^ b[14] ^ b[16] ^ b[17] ^ b[19] ^ b[21] ^ b[23] ^ b[24] ^ b[27] ^ b[28] ^ b[29] ^ b[33] ^ b[35] ^ b[37] ^ b[38] ^ b[39] ^ b[40] ^ b[43] ^ b[47] ^ b[49] ^ b[50] ^ b[51] ^ b[55] ^ b[57] ^ b[62];
	assign s[10] = p[10] ^ b[0] ^ b[1] ^ b[2] ^ b[3] ^ b[6] ^ b[7] ^ b[13] ^ b[14] ^ b[17] ^ b[18] ^ b[20] ^ b[22] ^ b[23] ^ b[24] ^ b[25] ^ b[27] ^ b[29] ^ b[30] ^ b[31] ^ b[32] ^ b[34] ^ b[35] ^ b[39] ^ b[43] ^ b[45] ^ b[46] ^ b[47] ^ b[49] ^ b[51] ^ b[58] ^ b[59] ^ b[63];

	assign en[0] = (s[4] ^ s[1]) | (s[5]) | (s[6] ^ s[1]) | (s[7] ^ s[0]) | (s[8] ^ s[0] ^ s[2] ^ s[3]) | (s[9] ^ s[0] ^ s[2]) | (s[10] ^ s[0] ^ s[1] ^ s[2] ^ s[3]);
	assign en[1] = (s[4] ^ s[1] ^ s[0]) | (s[5]) | (s[6] ^ s[1]) | (s[7]) | (s[8] ^ s[2] ^ s[3]) | (s[9] ^ s[2]) | (s[10] ^ s[1] ^ s[2] ^ s[3]);
	assign en[2] = (s[4] ^ s[0]) | (s[5] ^ s[1]) | (s[6] ^ s[1]) | (s[7] ^ s[1]) | (s[8] ^ s[2] ^ s[3] ^ s[1]) | (s[9] ^ s[2] ^ s[1]) | (s[10] ^ s[2] ^ s[3]);
	assign en[3] = (s[4] ^ s[0]) | (s[5] ^ s[1] ^ s[2]) | (s[6] ^ s[1]) | (s[7] ^ s[1] ^ s[2]) | (s[8] ^ s[3] ^ s[1]) | (s[9] ^ s[1] ^ s[2]) | (s[10] ^ s[3] ^ s[2]);
	assign en[4] = (s[4] ^ s[0]) | (s[5] ^ s[1] ^ s[2]) | (s[6] ^ s[1] ^ s[3]) | (s[7] ^ s[1] ^ s[2]) | (s[8] ^ s[1] ^ s[3]) | (s[9] ^ s[1] ^ s[2] ^ s[3]) | (s[10] ^ s[2] ^ s[3]);
	assign en[5] = (s[4] ^ s[0]) | (s[5] ^ s[1] ^ s[2] ^ s[0]) | (s[6] ^ s[1] ^ s[3]) | (s[7] ^ s[1] ^ s[2]) | (s[8] ^ s[1] ^ s[3] ^ s[0]) | (s[9] ^ s[1] ^ s[2] ^ s[3]) | (s[10] ^ s[2] ^ s[3]);
	assign en[6] = (s[4] ^ s[0]) | (s[5] ^ s[2] ^ s[0]) | (s[6] ^ s[3] ^ s[1]) | (s[7] ^ s[2] ^ s[1]) | (s[8] ^ s[3] ^ s[0] ^ s[1]) | (s[9] ^ s[2] ^ s[3]) | (s[10] ^ s[2] ^ s[3]);
	assign en[7] = (s[4] ^ s[0]) | (s[5] ^ s[0] ^ s[2]) | (s[6] ^ s[3] ^ s[1] ^ s[2]) | (s[7] ^ s[1]) | (s[8] ^ s[3] ^ s[0] ^ s[1]) | (s[9] ^ s[3]) | (s[10] ^ s[3]);
	assign en[8] = (s[4] ^ s[0]) | (s[5] ^ s[0] ^ s[2] ^ s[3]) | (s[6] ^ s[1] ^ s[2]) | (s[7] ^ s[1]) | (s[8] ^ s[0] ^ s[1]) | (s[9] ^ s[3]) | (s[10]);
	assign en[9] = (s[4]) | (s[5] ^ s[2] ^ s[3]) | (s[6] ^ s[1] ^ s[2]) | (s[7] ^ s[1] ^ s[0]) | (s[8] ^ s[1]) | (s[9] ^ s[3] ^ s[0]) | (s[10]);
	assign en[10] = (s[4]) | (s[5] ^ s[2] ^ s[3]) | (s[6] ^ s[2]) | (s[7] ^ s[0]) | (s[8]) | (s[9] ^ s[3] ^ s[0]) | (s[10] ^ s[1]);
	assign en[11] = (s[4]) | (s[5] ^ s[3] ^ s[2]) | (s[6] ^ s[2]) | (s[7] ^ s[0] ^ s[2]) | (s[8] ^ s[2]) | (s[9] ^ s[3] ^ s[0] ^ s[2]) | (s[10] ^ s[1] ^ s[2]);
	assign en[12] = (s[4] ^ s[3]) | (s[5] ^ s[2] ^ s[3]) | (s[6] ^ s[2] ^ s[3]) | (s[7] ^ s[0] ^ s[2] ^ s[3]) | (s[8] ^ s[2] ^ s[3]) | (s[9] ^ s[0] ^ s[2]) | (s[10] ^ s[1] ^ s[2]);
	assign en[13] = (s[4] ^ s[3] ^ s[0]) | (s[5] ^ s[2] ^ s[3] ^ s[0]) | (s[6] ^ s[2] ^ s[3]) | (s[7] ^ s[2] ^ s[3] ^ s[0]) | (s[8] ^ s[2] ^ s[3] ^ s[0]) | (s[9] ^ s[2] ^ s[0]) | (s[10] ^ s[1] ^ s[2]);
	assign en[14] = (s[4] ^ s[3] ^ s[0]) | (s[5] ^ s[2] ^ s[3] ^ s[0] ^ s[1]) | (s[6] ^ s[2] ^ s[3]) | (s[7] ^ s[2] ^ s[3] ^ s[0] ^ s[1]) | (s[8] ^ s[2] ^ s[3] ^ s[0] ^ s[1]) | (s[9] ^ s[2] ^ s[0] ^ s[1]) | (s[10] ^ s[2] ^ s[1]);
	assign en[15] = (s[4] ^ s[3] ^ s[0] ^ s[2]) | (s[5] ^ s[3] ^ s[0] ^ s[1]) | (s[6] ^ s[3] ^ s[2]) | (s[7] ^ s[3] ^ s[0] ^ s[1] ^ s[2]) | (s[8] ^ s[3] ^ s[0] ^ s[1]) | (s[9] ^ s[0] ^ s[1]) | (s[10] ^ s[1] ^ s[2]);
	assign en[16] = (s[4] ^ s[0] ^ s[2] ^ s[3]) | (s[5] ^ s[0] ^ s[1]) | (s[6] ^ s[2]) | (s[7] ^ s[0] ^ s[1] ^ s[2] ^ s[3]) | (s[8] ^ s[0] ^ s[1] ^ s[3]) | (s[9] ^ s[0] ^ s[1] ^ s[3]) | (s[10] ^ s[1] ^ s[2]);
	assign en[17] = (s[4] ^ s[2] ^ s[3]) | (s[5] ^ s[1] ^ s[0]) | (s[6] ^ s[2]) | (s[7] ^ s[1] ^ s[2] ^ s[3] ^ s[0]) | (s[8] ^ s[1] ^ s[3] ^ s[0]) | (s[9] ^ s[1] ^ s[3]) | (s[10] ^ s[1] ^ s[2] ^ s[0]);
	assign en[18] = (s[4] ^ s[2] ^ s[3]) | (s[5] ^ s[0]) | (s[6] ^ s[2] ^ s[1]) | (s[7] ^ s[2] ^ s[3] ^ s[0] ^ s[1]) | (s[8] ^ s[3] ^ s[0] ^ s[1]) | (s[9] ^ s[3] ^ s[1]) | (s[10] ^ s[2] ^ s[0]);
	assign en[19] = (s[4] ^ s[3] ^ s[2]) | (s[5] ^ s[0]) | (s[6] ^ s[1]) | (s[7] ^ s[3] ^ s[0] ^ s[1] ^ s[2]) | (s[8] ^ s[3] ^ s[0] ^ s[1]) | (s[9] ^ s[3] ^ s[1]) | (s[10] ^ s[0] ^ s[2]);
	assign en[20] = (s[4] ^ s[2]) | (s[5] ^ s[0]) | (s[6] ^ s[1] ^ s[3]) | (s[7] ^ s[0] ^ s[1] ^ s[2]) | (s[8] ^ s[0] ^ s[1]) | (s[9] ^ s[1] ^ s[3]) | (s[10] ^ s[0] ^ s[2] ^ s[3]);
	assign en[21] = (s[4] ^ s[2]) | (s[5]) | (s[6] ^ s[1] ^ s[3]) | (s[7] ^ s[1] ^ s[2] ^ s[0]) | (s[8] ^ s[1]) | (s[9] ^ s[1] ^ s[3] ^ s[0]) | (s[10] ^ s[2] ^ s[3] ^ s[0]);
	assign en[22] = (s[4] ^ s[2] ^ s[1]) | (s[5]) | (s[6] ^ s[3]) | (s[7] ^ s[2] ^ s[0]) | (s[8]) | (s[9] ^ s[3] ^ s[0]) | (s[10] ^ s[2] ^ s[3] ^ s[0] ^ s[1]);
	assign en[23] = (s[4] ^ s[1]) | (s[5] ^ s[2]) | (s[6] ^ s[3]) | (s[7] ^ s[0] ^ s[2]) | (s[8]) | (s[9] ^ s[3] ^ s[0]) | (s[10] ^ s[3] ^ s[0] ^ s[1]);
	assign en[24] = (s[4] ^ s[1]) | (s[5] ^ s[2]) | (s[6]) | (s[7] ^ s[0] ^ s[2]) | (s[8]) | (s[9] ^ s[0] ^ s[3]) | (s[10] ^ s[0] ^ s[1] ^ s[3]);
	assign en[25] = (s[4] ^ s[1] ^ s[0]) | (s[5] ^ s[2] ^ s[0]) | (s[6] ^ s[0]) | (s[7] ^ s[2] ^ s[0]) | (s[8] ^ s[0]) | (s[9] ^ s[3] ^ s[0]) | (s[10] ^ s[1] ^ s[3]);
	assign en[26] = (s[4] ^ s[0] ^ s[1]) | (s[5] ^ s[2] ^ s[0]) | (s[6] ^ s[0] ^ s[1]) | (s[7] ^ s[2] ^ s[0] ^ s[1]) | (s[8] ^ s[0] ^ s[1]) | (s[9] ^ s[3] ^ s[0] ^ s[1]) | (s[10] ^ s[3] ^ s[1]);
	assign en[27] = (s[4] ^ s[0] ^ s[1] ^ s[2]) | (s[5] ^ s[0] ^ s[2]) | (s[6] ^ s[0] ^ s[1] ^ s[2]) | (s[7] ^ s[0] ^ s[1] ^ s[2]) | (s[8] ^ s[0] ^ s[1]) | (s[9] ^ s[3] ^ s[0] ^ s[1]) | (s[10] ^ s[3] ^ s[1] ^ s[2]);
	assign en[28] = (s[4] ^ s[0] ^ s[1] ^ s[2] ^ s[3]) | (s[5] ^ s[0] ^ s[2]) | (s[6] ^ s[0] ^ s[1] ^ s[2] ^ s[3]) | (s[7] ^ s[0] ^ s[1] ^ s[2] ^ s[3]) | (s[8] ^ s[0] ^ s[1] ^ s[3]) | (s[9] ^ s[0] ^ s[1]) | (s[10] ^ s[1] ^ s[2] ^ s[3]);
	assign en[29] = (s[4] ^ s[1] ^ s[2] ^ s[3]) | (s[5] ^ s[2] ^ s[0]) | (s[6] ^ s[1] ^ s[2] ^ s[3] ^ s[0]) | (s[7] ^ s[1] ^ s[2] ^ s[3] ^ s[0]) | (s[8] ^ s[1] ^ s[3] ^ s[0]) | (s[9] ^ s[1]) | (s[10] ^ s[1] ^ s[2] ^ s[3] ^ s[0]);
	assign en[30] = (s[4] ^ s[2] ^ s[3] ^ s[1]) | (s[5] ^ s[2] ^ s[0] ^ s[1]) | (s[6] ^ s[2] ^ s[3] ^ s[0]) | (s[7] ^ s[2] ^ s[3] ^ s[0] ^ s[1]) | (s[8] ^ s[3] ^ s[0]) | (s[9] ^ s[1]) | (s[10] ^ s[2] ^ s[3] ^ s[0]);
	assign en[31] = (s[4] ^ s[3] ^ s[1] ^ s[2]) | (s[5] ^ s[0] ^ s[1] ^ s[2]) | (s[6] ^ s[3] ^ s[0]) | (s[7] ^ s[3] ^ s[0] ^ s[1]) | (s[8] ^ s[3] ^ s[0] ^ s[2]) | (s[9] ^ s[1]) | (s[10] ^ s[3] ^ s[0] ^ s[2]);
	assign en[32] = (s[4] ^ s[1] ^ s[2] ^ s[3]) | (s[5] ^ s[0] ^ s[1] ^ s[2]) | (s[6] ^ s[0]) | (s[7] ^ s[0] ^ s[1]) | (s[8] ^ s[0] ^ s[2] ^ s[3]) | (s[9] ^ s[1] ^ s[3]) | (s[10] ^ s[0] ^ s[2] ^ s[3]);
	assign en[33] = (s[4] ^ s[1] ^ s[2] ^ s[3]) | (s[5] ^ s[1] ^ s[2] ^ s[0]) | (s[6] ^ s[0]) | (s[7] ^ s[1] ^ s[0]) | (s[8] ^ s[2] ^ s[3] ^ s[0]) | (s[9] ^ s[1] ^ s[3]) | (s[10] ^ s[2] ^ s[3]);
	assign en[34] = (s[4] ^ s[2] ^ s[3]) | (s[5] ^ s[2] ^ s[0] ^ s[1]) | (s[6] ^ s[0]) | (s[7] ^ s[0] ^ s[1]) | (s[8] ^ s[2] ^ s[3] ^ s[0] ^ s[1]) | (s[9] ^ s[3] ^ s[1]) | (s[10] ^ s[2] ^ s[3]);
	assign en[35] = (s[4] ^ s[3]) | (s[5] ^ s[0] ^ s[1]) | (s[6] ^ s[0] ^ s[2]) | (s[7] ^ s[0] ^ s[1] ^ s[2]) | (s[8] ^ s[3] ^ s[0] ^ s[1] ^ s[2]) | (s[9] ^ s[3] ^ s[1] ^ s[2]) | (s[10] ^ s[3]);
	assign en[36] = (s[4]) | (s[5] ^ s[0] ^ s[1]) | (s[6] ^ s[0] ^ s[2] ^ s[3]) | (s[7] ^ s[0] ^ s[1] ^ s[2] ^ s[3]) | (s[8] ^ s[0] ^ s[1] ^ s[2]) | (s[9] ^ s[1] ^ s[2] ^ s[3]) | (s[10] ^ s[3]);
	assign en[37] = (s[4] ^ s[0]) | (s[5] ^ s[1] ^ s[0]) | (s[6] ^ s[2] ^ s[3]) | (s[7] ^ s[1] ^ s[2] ^ s[3]) | (s[8] ^ s[1] ^ s[2]) | (s[9] ^ s[1] ^ s[2] ^ s[3] ^ s[0]) | (s[10] ^ s[3]);
	assign en[38] = (s[4] ^ s[0] ^ s[1]) | (s[5] ^ s[0]) | (s[6] ^ s[2] ^ s[3] ^ s[1]) | (s[7] ^ s[2] ^ s[3] ^ s[1]) | (s[8] ^ s[2]) | (s[9] ^ s[2] ^ s[3] ^ s[0]) | (s[10] ^ s[3]);
	assign en[39] = (s[4] ^ s[0] ^ s[1] ^ s[2]) | (s[5] ^ s[0]) | (s[6] ^ s[3] ^ s[1]) | (s[7] ^ s[3] ^ s[1] ^ s[2]) | (s[8] ^ s[2]) | (s[9] ^ s[3] ^ s[0]) | (s[10] ^ s[3]);
	assign en[40] = (s[4] ^ s[0] ^ s[1] ^ s[2] ^ s[3]) | (s[5] ^ s[0]) | (s[6] ^ s[1]) | (s[7] ^ s[1] ^ s[2]) | (s[8] ^ s[2]) | (s[9] ^ s[0] ^ s[3]) | (s[10] ^ s[3]);
	assign en[41] = (s[4] ^ s[1] ^ s[2] ^ s[3]) | (s[5] ^ s[0]) | (s[6] ^ s[1] ^ s[0]) | (s[7] ^ s[1] ^ s[2]) | (s[8] ^ s[2] ^ s[0]) | (s[9] ^ s[3]) | (s[10] ^ s[3]);
	assign en[42] = (s[4] ^ s[2] ^ s[3]) | (s[5] ^ s[0] ^ s[1]) | (s[6] ^ s[0]) | (s[7] ^ s[2] ^ s[1]) | (s[8] ^ s[2] ^ s[0]) | (s[9] ^ s[3]) | (s[10] ^ s[3] ^ s[1]);
	assign en[43] = (s[4] ^ s[3]) | (s[5] ^ s[0] ^ s[1] ^ s[2]) | (s[6] ^ s[0]) | (s[7] ^ s[1]) | (s[8] ^ s[0] ^ s[2]) | (s[9] ^ s[3]) | (s[10] ^ s[3] ^ s[1] ^ s[2]);
	assign en[44] = (s[4]) | (s[5] ^ s[0] ^ s[1] ^ s[2] ^ s[3]) | (s[6] ^ s[0]) | (s[7] ^ s[1]) | (s[8] ^ s[0] ^ s[2]) | (s[9] ^ s[3]) | (s[10] ^ s[1] ^ s[2] ^ s[3]);
	assign en[45] = (s[4]) | (s[5] ^ s[1] ^ s[2] ^ s[3]) | (s[6] ^ s[0]) | (s[7] ^ s[1] ^ s[0]) | (s[8] ^ s[2] ^ s[0]) | (s[9] ^ s[3]) | (s[10] ^ s[1] ^ s[2] ^ s[3]);
	assign en[46] = (s[4]) | (s[5] ^ s[2] ^ s[3]) | (s[6] ^ s[0] ^ s[1]) | (s[7] ^ s[0]) | (s[8] ^ s[2] ^ s[0]) | (s[9] ^ s[3] ^ s[1]) | (s[10] ^ s[2] ^ s[3] ^ s[1]);
	assign en[47] = (s[4]) | (s[5] ^ s[3]) | (s[6] ^ s[0] ^ s[1]) | (s[7] ^ s[0] ^ s[2]) | (s[8] ^ s[0] ^ s[2]) | (s[9] ^ s[3] ^ s[1] ^ s[2]) | (s[10] ^ s[3] ^ s[1]);
	assign en[48] = (s[4]) | (s[5]) | (s[6] ^ s[0] ^ s[1]) | (s[7] ^ s[0] ^ s[2]) | (s[8] ^ s[0] ^ s[2] ^ s[3]) | (s[9] ^ s[1] ^ s[2] ^ s[3]) | (s[10] ^ s[1] ^ s[3]);
	assign en[49] = (s[4] ^ s[0]) | (s[5] ^ s[0]) | (s[6] ^ s[1]) | (s[7] ^ s[2]) | (s[8] ^ s[2] ^ s[3]) | (s[9] ^ s[1] ^ s[2] ^ s[3]) | (s[10] ^ s[1] ^ s[3]);
	assign en[50] = (s[4] ^ s[0] ^ s[1]) | (s[5] ^ s[0]) | (s[6] ^ s[1]) | (s[7] ^ s[2]) | (s[8] ^ s[2] ^ s[3]) | (s[9] ^ s[2] ^ s[3]) | (s[10] ^ s[3]);
	assign en[51] = (s[4] ^ s[0] ^ s[1] ^ s[2]) | (s[5] ^ s[0]) | (s[6] ^ s[1]) | (s[7] ^ s[2]) | (s[8] ^ s[3]) | (s[9] ^ s[3]) | (s[10] ^ s[3]);
	assign en[52] = (s[4] ^ s[0] ^ s[1] ^ s[2] ^ s[3]) | (s[5] ^ s[0]) | (s[6] ^ s[1]) | (s[7] ^ s[2]) | (s[8]) | (s[9] ^ s[3]) | (s[10]);
	assign en[53] = (s[4] ^ s[1] ^ s[2] ^ s[3]) | (s[5] ^ s[0]) | (s[6] ^ s[1]) | (s[7] ^ s[2]) | (s[8] ^ s[0]) | (s[9] ^ s[3]) | (s[10]);
	assign en[54] = (s[4] ^ s[2] ^ s[3]) | (s[5] ^ s[0] ^ s[1]) | (s[6]) | (s[7] ^ s[2]) | (s[8] ^ s[0]) | (s[9] ^ s[3] ^ s[1]) | (s[10]);
	assign en[55] = (s[4] ^ s[3]) | (s[5] ^ s[0] ^ s[1] ^ s[2]) | (s[6]) | (s[7]) | (s[8] ^ s[0]) | (s[9] ^ s[3] ^ s[1]) | (s[10] ^ s[2]);
	assign en[56] = (s[4]) | (s[5] ^ s[0] ^ s[1] ^ s[2]) | (s[6] ^ s[3]) | (s[7]) | (s[8] ^ s[0]) | (s[9] ^ s[1]) | (s[10] ^ s[2] ^ s[3]);
	assign en[57] = (s[4]) | (s[5] ^ s[1] ^ s[2]) | (s[6] ^ s[3]) | (s[7] ^ s[0]) | (s[8]) | (s[9] ^ s[1]) | (s[10] ^ s[2] ^ s[3]);
	assign en[58] = (s[4]) | (s[5] ^ s[2]) | (s[6] ^ s[3]) | (s[7] ^ s[0]) | (s[8] ^ s[1]) | (s[9]) | (s[10] ^ s[2] ^ s[3]);
	assign en[59] = (s[4]) | (s[5]) | (s[6] ^ s[3]) | (s[7] ^ s[0]) | (s[8] ^ s[1]) | (s[9] ^ s[2]) | (s[10] ^ s[3]);
	assign en[60] = (s[4]) | (s[5]) | (s[6]) | (s[7] ^ s[0]) | (s[8] ^ s[1]) | (s[9] ^ s[2]) | (s[10] ^ s[3]);
	assign en[61] = (s[4]) | (s[5]) | (s[6]) | (s[7]) | (s[8] ^ s[1]) | (s[9] ^ s[2]) | (s[10] ^ s[3]);
	assign en[62] = (s[4]) | (s[5]) | (s[6]) | (s[7]) | (s[8]) | (s[9] ^ s[2]) | (s[10] ^ s[3]);
	assign en[63] = (s[4]) | (s[5]) | (s[6]) | (s[7]) | (s[8]) | (s[9]) | (s[10] ^ s[3]);

	assign m[0] = ((~( en[0] )) & s[0]) ^ b[0];
	assign m[1] = ((~( en[1] & en[0] )) & s[1]) ^ b[1];
	assign m[2] = ((~( en[2] & en[1] & en[0] )) & s[2]) ^ b[2];
	assign m[3] = ((~( en[3] & en[2] & en[1] & en[0] )) & s[3]) ^ b[3];
	assign m[4] = ((~( en[4] & en[3] & en[2] & en[1] )) & s[0]) ^ b[4];
	assign m[5] = ((~( en[5] & en[4] & en[3] & en[2] )) & s[1]) ^ b[5];
	assign m[6] = ((~( en[6] & en[5] & en[4] & en[3] )) & s[2]) ^ b[6];
	assign m[7] = ((~( en[7] & en[6] & en[5] & en[4] )) & s[3]) ^ b[7];
	assign m[8] = ((~( en[8] & en[7] & en[6] & en[5] )) & s[0]) ^ b[8];
	assign m[9] = ((~( en[9] & en[8] & en[7] & en[6] )) & s[1]) ^ b[9];
	assign m[10] = ((~( en[10] & en[9] & en[8] & en[7] )) & s[2]) ^ b[10];
	assign m[11] = ((~( en[11] & en[10] & en[9] & en[8] )) & s[3]) ^ b[11];
	assign m[12] = ((~( en[12] & en[11] & en[10] & en[9] )) & s[0]) ^ b[12];
	assign m[13] = ((~( en[13] & en[12] & en[11] & en[10] )) & s[1]) ^ b[13];
	assign m[14] = ((~( en[14] & en[13] & en[12] & en[11] )) & s[2]) ^ b[14];
	assign m[15] = ((~( en[15] & en[14] & en[13] & en[12] )) & s[3]) ^ b[15];
	assign m[16] = ((~( en[16] & en[15] & en[14] & en[13] )) & s[0]) ^ b[16];
	assign m[17] = ((~( en[17] & en[16] & en[15] & en[14] )) & s[1]) ^ b[17];
	assign m[18] = ((~( en[18] & en[17] & en[16] & en[15] )) & s[2]) ^ b[18];
	assign m[19] = ((~( en[19] & en[18] & en[17] & en[16] )) & s[3]) ^ b[19];
	assign m[20] = ((~( en[20] & en[19] & en[18] & en[17] )) & s[0]) ^ b[20];
	assign m[21] = ((~( en[21] & en[20] & en[19] & en[18] )) & s[1]) ^ b[21];
	assign m[22] = ((~( en[22] & en[21] & en[20] & en[19] )) & s[2]) ^ b[22];
	assign m[23] = ((~( en[23] & en[22] & en[21] & en[20] )) & s[3]) ^ b[23];
	assign m[24] = ((~( en[24] & en[23] & en[22] & en[21] )) & s[0]) ^ b[24];
	assign m[25] = ((~( en[25] & en[24] & en[23] & en[22] )) & s[1]) ^ b[25];
	assign m[26] = ((~( en[26] & en[25] & en[24] & en[23] )) & s[2]) ^ b[26];
	assign m[27] = ((~( en[27] & en[26] & en[25] & en[24] )) & s[3]) ^ b[27];
	assign m[28] = ((~( en[28] & en[27] & en[26] & en[25] )) & s[0]) ^ b[28];
	assign m[29] = ((~( en[29] & en[28] & en[27] & en[26] )) & s[1]) ^ b[29];
	assign m[30] = ((~( en[30] & en[29] & en[28] & en[27] )) & s[2]) ^ b[30];
	assign m[31] = ((~( en[31] & en[30] & en[29] & en[28] )) & s[3]) ^ b[31];
	assign m[32] = ((~( en[32] & en[31] & en[30] & en[29] )) & s[0]) ^ b[32];
	assign m[33] = ((~( en[33] & en[32] & en[31] & en[30] )) & s[1]) ^ b[33];
	assign m[34] = ((~( en[34] & en[33] & en[32] & en[31] )) & s[2]) ^ b[34];
	assign m[35] = ((~( en[35] & en[34] & en[33] & en[32] )) & s[3]) ^ b[35];
	assign m[36] = ((~( en[36] & en[35] & en[34] & en[33] )) & s[0]) ^ b[36];
	assign m[37] = ((~( en[37] & en[36] & en[35] & en[34] )) & s[1]) ^ b[37];
	assign m[38] = ((~( en[38] & en[37] & en[36] & en[35] )) & s[2]) ^ b[38];
	assign m[39] = ((~( en[39] & en[38] & en[37] & en[36] )) & s[3]) ^ b[39];
	assign m[40] = ((~( en[40] & en[39] & en[38] & en[37] )) & s[0]) ^ b[40];
	assign m[41] = ((~( en[41] & en[40] & en[39] & en[38] )) & s[1]) ^ b[41];
	assign m[42] = ((~( en[42] & en[41] & en[40] & en[39] )) & s[2]) ^ b[42];
	assign m[43] = ((~( en[43] & en[42] & en[41] & en[40] )) & s[3]) ^ b[43];
	assign m[44] = ((~( en[44] & en[43] & en[42] & en[41] )) & s[0]) ^ b[44];
	assign m[45] = ((~( en[45] & en[44] & en[43] & en[42] )) & s[1]) ^ b[45];
	assign m[46] = ((~( en[46] & en[45] & en[44] & en[43] )) & s[2]) ^ b[46];
	assign m[47] = ((~( en[47] & en[46] & en[45] & en[44] )) & s[3]) ^ b[47];
	assign m[48] = ((~( en[48] & en[47] & en[46] & en[45] )) & s[0]) ^ b[48];
	assign m[49] = ((~( en[49] & en[48] & en[47] & en[46] )) & s[1]) ^ b[49];
	assign m[50] = ((~( en[50] & en[49] & en[48] & en[47] )) & s[2]) ^ b[50];
	assign m[51] = ((~( en[51] & en[50] & en[49] & en[48] )) & s[3]) ^ b[51];
	assign m[52] = ((~( en[52] & en[51] & en[50] & en[49] )) & s[0]) ^ b[52];
	assign m[53] = ((~( en[53] & en[52] & en[51] & en[50] )) & s[1]) ^ b[53];
	assign m[54] = ((~( en[54] & en[53] & en[52] & en[51] )) & s[2]) ^ b[54];
	assign m[55] = ((~( en[55] & en[54] & en[53] & en[52] )) & s[3]) ^ b[55];
	assign m[56] = ((~( en[56] & en[55] & en[54] & en[53] )) & s[0]) ^ b[56];
	assign m[57] = ((~( en[57] & en[56] & en[55] & en[54] )) & s[1]) ^ b[57];
	assign m[58] = ((~( en[58] & en[57] & en[56] & en[55] )) & s[2]) ^ b[58];
	assign m[59] = ((~( en[59] & en[58] & en[57] & en[56] )) & s[3]) ^ b[59];
	assign m[60] = ((~( en[60] & en[59] & en[58] & en[57] )) & s[0]) ^ b[60];
	assign m[61] = ((~( en[61] & en[60] & en[59] & en[58] )) & s[1]) ^ b[61];
	assign m[62] = ((~( en[62] & en[61] & en[60] & en[59] )) & s[2]) ^ b[62];
	assign m[63] = ((~( en[63] & en[62] & en[61] & en[60] )) & s[3]) ^ b[63];

endmodule