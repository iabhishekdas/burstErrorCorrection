module encoder (
	input [0:31] m,
	output [0:40] c
);

	wire [0:8] p;

	assign p[0] = m[2] ^ m[5] ^ m[8] ^ m[11] ^ m[14] ^ m[17] ^ m[20] ^ m[23] ^ m[26] ^ m[29] ^ 0;
	assign p[1] = m[0] ^ m[3] ^ m[6] ^ m[9] ^ m[12] ^ m[15] ^ m[18] ^ m[21] ^ m[24] ^ m[27] ^ m[30] ^ 0;
	assign p[2] = m[1] ^ m[4] ^ m[7] ^ m[10] ^ m[13] ^ m[16] ^ m[19] ^ m[22] ^ m[25] ^ m[28] ^ m[31] ^ 0;
	assign p[3] = m[0] ^ m[4] ^ m[5] ^ m[6] ^ m[7] ^ m[10] ^ m[11] ^ m[12] ^ m[16] ^ m[17] ^ m[26] ^ 0;
	assign p[4] = m[4] ^ m[5] ^ m[8] ^ m[10] ^ m[13] ^ m[14] ^ m[18] ^ m[19] ^ m[20] ^ m[21] ^ m[27] ^ 0;
	assign p[5] = m[2] ^ m[6] ^ m[8] ^ m[9] ^ m[13] ^ m[15] ^ m[16] ^ m[18] ^ m[22] ^ m[23] ^ m[28] ^ 0;
	assign p[6] = m[0] ^ m[1] ^ m[4] ^ m[6] ^ m[7] ^ m[8] ^ m[9] ^ m[11] ^ m[14] ^ m[19] ^ m[24] ^ m[29] ^ 0;
	assign p[7] = m[4] ^ m[5] ^ m[6] ^ m[7] ^ m[9] ^ m[11] ^ m[12] ^ m[13] ^ m[15] ^ m[20] ^ m[22] ^ m[25] ^ m[30] ^ 0;
	assign p[8] = m[1] ^ m[3] ^ m[4] ^ m[5] ^ m[7] ^ m[8] ^ m[9] ^ m[10] ^ m[12] ^ m[14] ^ m[15] ^ m[17] ^ m[21] ^ m[23] ^ m[24] ^ m[25] ^ m[31] ^ 0;

	assign c = {m,p};

endmodule

module decoder (
	input [0:40] c,
	output [0:31] m
);

	wire [0:8] p, s;
	wire [0:31] b, en;
	assign b = c[0:31];
	assign p = c[32:40];

	assign s[0] = p[0] ^ b[2] ^ b[5] ^ b[8] ^ b[11] ^ b[14] ^ b[17] ^ b[20] ^ b[23] ^ b[26] ^ b[29] ^ 0;
	assign s[1] = p[1] ^ b[0] ^ b[3] ^ b[6] ^ b[9] ^ b[12] ^ b[15] ^ b[18] ^ b[21] ^ b[24] ^ b[27] ^ b[30] ^ 0;
	assign s[2] = p[2] ^ b[1] ^ b[4] ^ b[7] ^ b[10] ^ b[13] ^ b[16] ^ b[19] ^ b[22] ^ b[25] ^ b[28] ^ b[31] ^ 0;
	assign s[3] = p[3] ^ b[0] ^ b[4] ^ b[5] ^ b[6] ^ b[7] ^ b[10] ^ b[11] ^ b[12] ^ b[16] ^ b[17] ^ b[26] ^ 0;
	assign s[4] = p[4] ^ b[4] ^ b[5] ^ b[8] ^ b[10] ^ b[13] ^ b[14] ^ b[18] ^ b[19] ^ b[20] ^ b[21] ^ b[27] ^ 0;
	assign s[5] = p[5] ^ b[2] ^ b[6] ^ b[8] ^ b[9] ^ b[13] ^ b[15] ^ b[16] ^ b[18] ^ b[22] ^ b[23] ^ b[28] ^ 0;
	assign s[6] = p[6] ^ b[0] ^ b[1] ^ b[4] ^ b[6] ^ b[7] ^ b[8] ^ b[9] ^ b[11] ^ b[14] ^ b[19] ^ b[24] ^ b[29] ^ 0;
	assign s[7] = p[7] ^ b[4] ^ b[5] ^ b[6] ^ b[7] ^ b[9] ^ b[11] ^ b[12] ^ b[13] ^ b[15] ^ b[20] ^ b[22] ^ b[25] ^ b[30] ^ 0;
	assign s[8] = p[8] ^ b[1] ^ b[3] ^ b[4] ^ b[5] ^ b[7] ^ b[8] ^ b[9] ^ b[10] ^ b[12] ^ b[14] ^ b[15] ^ b[17] ^ b[21] ^ b[23] ^ b[24] ^ b[25] ^ b[31] ^ 0;

	assign en[0] = (s[3] ^ s[1] ^ 0) | (s[4] ^ 0) | (s[5] ^ s[0] ^ 0) | (s[6] ^ s[1] ^ s[2] ^ 0) | (s[7] ^ 0) | (s[8] ^ s[2] ^ 0);
	assign en[1] = (s[3] ^ 0) | (s[4] ^ 0) | (s[5] ^ s[0] ^ 0) | (s[6] ^ s[2] ^ 0) | (s[7] ^ 0) | (s[8] ^ s[2] ^ s[1] ^ 0);
	assign en[2] = (s[3] ^ s[2] ^ 0) | (s[4] ^ s[2] ^ 0) | (s[5] ^ s[0] ^ 0) | (s[6] ^ s[2] ^ 0) | (s[7] ^ s[2] ^ 0) | (s[8] ^ s[1] ^ s[2] ^ 0);
	assign en[3] = (s[3] ^ s[2] ^ s[0] ^ 0) | (s[4] ^ s[2] ^ s[0] ^ 0) | (s[5] ^ 0) | (s[6] ^ s[2] ^ 0) | (s[7] ^ s[2] ^ s[0] ^ 0) | (s[8] ^ s[1] ^ s[2] ^ s[0] ^ 0);
	assign en[4] = (s[3] ^ s[2] ^ s[0] ^ s[1] ^ 0) | (s[4] ^ s[2] ^ s[0] ^ 0) | (s[5] ^ s[1] ^ 0) | (s[6] ^ s[2] ^ s[1] ^ 0) | (s[7] ^ s[2] ^ s[0] ^ s[1] ^ 0) | (s[8] ^ s[2] ^ s[0] ^ 0);
	assign en[5] = (s[3] ^ s[0] ^ s[1] ^ s[2] ^ 0) | (s[4] ^ s[0] ^ 0) | (s[5] ^ s[1] ^ 0) | (s[6] ^ s[1] ^ s[2] ^ 0) | (s[7] ^ s[0] ^ s[1] ^ s[2] ^ 0) | (s[8] ^ s[0] ^ s[2] ^ 0);
	assign en[6] = (s[3] ^ s[1] ^ s[2] ^ 0) | (s[4] ^ s[0] ^ 0) | (s[5] ^ s[1] ^ s[0] ^ 0) | (s[6] ^ s[1] ^ s[2] ^ s[0] ^ 0) | (s[7] ^ s[1] ^ s[2] ^ 0) | (s[8] ^ s[2] ^ s[0] ^ 0);
	assign en[7] = (s[3] ^ s[2] ^ 0) | (s[4] ^ s[0] ^ 0) | (s[5] ^ s[0] ^ s[1] ^ 0) | (s[6] ^ s[2] ^ s[0] ^ s[1] ^ 0) | (s[7] ^ s[2] ^ s[1] ^ 0) | (s[8] ^ s[2] ^ s[0] ^ s[1] ^ 0);
	assign en[8] = (s[3] ^ s[2] ^ 0) | (s[4] ^ s[0] ^ s[2] ^ 0) | (s[5] ^ s[0] ^ s[1] ^ 0) | (s[6] ^ s[0] ^ s[1] ^ 0) | (s[7] ^ s[1] ^ 0) | (s[8] ^ s[0] ^ s[1] ^ s[2] ^ 0);
	assign en[9] = (s[3] ^ s[2] ^ s[0] ^ 0) | (s[4] ^ s[2] ^ 0) | (s[5] ^ s[1] ^ 0) | (s[6] ^ s[1] ^ s[0] ^ 0) | (s[7] ^ s[1] ^ s[0] ^ 0) | (s[8] ^ s[1] ^ s[2] ^ 0);
	assign en[10] = (s[3] ^ s[2] ^ s[0] ^ s[1] ^ 0) | (s[4] ^ s[2] ^ 0) | (s[5] ^ 0) | (s[6] ^ s[0] ^ 0) | (s[7] ^ s[0] ^ s[1] ^ 0) | (s[8] ^ s[2] ^ s[1] ^ 0);
	assign en[11] = (s[3] ^ s[0] ^ s[1] ^ 0) | (s[4] ^ s[2] ^ 0) | (s[5] ^ s[2] ^ 0) | (s[6] ^ s[0] ^ 0) | (s[7] ^ s[0] ^ s[1] ^ s[2] ^ 0) | (s[8] ^ s[1] ^ 0);
	assign en[12] = (s[3] ^ s[1] ^ 0) | (s[4] ^ s[2] ^ s[0] ^ 0) | (s[5] ^ s[2] ^ 0) | (s[6] ^ s[0] ^ 0) | (s[7] ^ s[1] ^ s[2] ^ 0) | (s[8] ^ s[1] ^ s[0] ^ 0);
	assign en[13] = (s[3] ^ 0) | (s[4] ^ s[2] ^ s[0] ^ 0) | (s[5] ^ s[2] ^ s[1] ^ 0) | (s[6] ^ s[0] ^ 0) | (s[7] ^ s[2] ^ s[1] ^ 0) | (s[8] ^ s[0] ^ s[1] ^ 0);
	assign en[14] = (s[3] ^ s[2] ^ 0) | (s[4] ^ s[0] ^ 0) | (s[5] ^ s[1] ^ s[2] ^ 0) | (s[6] ^ s[0] ^ 0) | (s[7] ^ s[1] ^ 0) | (s[8] ^ s[0] ^ s[1] ^ 0);
	assign en[15] = (s[3] ^ s[2] ^ s[0] ^ 0) | (s[4] ^ 0) | (s[5] ^ s[1] ^ s[2] ^ 0) | (s[6] ^ 0) | (s[7] ^ s[1] ^ 0) | (s[8] ^ s[1] ^ s[0] ^ 0);
	assign en[16] = (s[3] ^ s[2] ^ s[0] ^ 0) | (s[4] ^ s[1] ^ 0) | (s[5] ^ s[2] ^ s[1] ^ 0) | (s[6] ^ 0) | (s[7] ^ 0) | (s[8] ^ s[0] ^ 0);
	assign en[17] = (s[3] ^ s[0] ^ 0) | (s[4] ^ s[1] ^ s[2] ^ 0) | (s[5] ^ s[1] ^ 0) | (s[6] ^ s[2] ^ 0) | (s[7] ^ 0) | (s[8] ^ s[0] ^ 0);
	assign en[18] = (s[3] ^ 0) | (s[4] ^ s[1] ^ s[2] ^ s[0] ^ 0) | (s[5] ^ s[1] ^ 0) | (s[6] ^ s[2] ^ 0) | (s[7] ^ s[0] ^ 0) | (s[8] ^ 0);
	assign en[19] = (s[3] ^ 0) | (s[4] ^ s[2] ^ s[0] ^ s[1] ^ 0) | (s[5] ^ 0) | (s[6] ^ s[2] ^ 0) | (s[7] ^ s[0] ^ 0) | (s[8] ^ s[1] ^ 0);
	assign en[20] = (s[3] ^ 0) | (s[4] ^ s[0] ^ s[1] ^ 0) | (s[5] ^ s[2] ^ 0) | (s[6] ^ 0) | (s[7] ^ s[0] ^ s[2] ^ 0) | (s[8] ^ s[1] ^ 0);
	assign en[21] = (s[3] ^ 0) | (s[4] ^ s[1] ^ 0) | (s[5] ^ s[2] ^ s[0] ^ 0) | (s[6] ^ 0) | (s[7] ^ s[2] ^ 0) | (s[8] ^ s[1] ^ s[0] ^ 0);
	assign en[22] = (s[3] ^ 0) | (s[4] ^ 0) | (s[5] ^ s[2] ^ s[0] ^ 0) | (s[6] ^ s[1] ^ 0) | (s[7] ^ s[2] ^ 0) | (s[8] ^ s[0] ^ s[1] ^ 0);
	assign en[23] = (s[3] ^ 0) | (s[4] ^ 0) | (s[5] ^ s[0] ^ 0) | (s[6] ^ s[1] ^ 0) | (s[7] ^ s[2] ^ 0) | (s[8] ^ s[0] ^ s[1] ^ s[2] ^ 0);
	assign en[24] = (s[3] ^ s[0] ^ 0) | (s[4] ^ 0) | (s[5] ^ 0) | (s[6] ^ s[1] ^ 0) | (s[7] ^ s[2] ^ 0) | (s[8] ^ s[1] ^ s[2] ^ 0);
	assign en[25] = (s[3] ^ s[0] ^ 0) | (s[4] ^ s[1] ^ 0) | (s[5] ^ 0) | (s[6] ^ 0) | (s[7] ^ s[2] ^ 0) | (s[8] ^ s[2] ^ 0);
	assign en[26] = (s[3] ^ s[0] ^ 0) | (s[4] ^ s[1] ^ 0) | (s[5] ^ s[2] ^ 0) | (s[6] ^ 0) | (s[7] ^ 0) | (s[8] ^ 0);
	assign en[27] = (s[3] ^ 0) | (s[4] ^ s[1] ^ 0) | (s[5] ^ s[2] ^ 0) | (s[6] ^ s[0] ^ 0) | (s[7] ^ 0) | (s[8] ^ 0);
	assign en[28] = (s[3] ^ 0) | (s[4] ^ 0) | (s[5] ^ s[2] ^ 0) | (s[6] ^ s[0] ^ 0) | (s[7] ^ s[1] ^ 0) | (s[8] ^ 0);
	assign en[29] = (s[3] ^ 0) | (s[4] ^ 0) | (s[5] ^ 0) | (s[6] ^ s[0] ^ 0) | (s[7] ^ s[1] ^ 0) | (s[8] ^ s[2] ^ 0);
	assign en[30] = (s[3] ^ 0) | (s[4] ^ 0) | (s[5] ^ 0) | (s[6] ^ 0) | (s[7] ^ s[1] ^ 0) | (s[8] ^ s[2] ^ 0);
	assign en[31] = (s[3] ^ 0) | (s[4] ^ 0) | (s[5] ^ 0) | (s[6] ^ 0) | (s[7] ^ 0) | (s[8] ^ s[2] ^ 0);

	assign m[0] = ((~( en[0] )) & s[1]) ^ b[0];
	assign m[1] = ((~( en[1] & en[0] )) & s[2]) ^ b[1];
	assign m[2] = ((~( en[2] & en[1] & en[0] )) & s[0]) ^ b[2];
	assign m[3] = ((~( en[3] & en[2] & en[1] )) & s[1]) ^ b[3];
	assign m[4] = ((~( en[4] & en[3] & en[2] )) & s[2]) ^ b[4];
	assign m[5] = ((~( en[5] & en[4] & en[3] )) & s[0]) ^ b[5];
	assign m[6] = ((~( en[6] & en[5] & en[4] )) & s[1]) ^ b[6];
	assign m[7] = ((~( en[7] & en[6] & en[5] )) & s[2]) ^ b[7];
	assign m[8] = ((~( en[8] & en[7] & en[6] )) & s[0]) ^ b[8];
	assign m[9] = ((~( en[9] & en[8] & en[7] )) & s[1]) ^ b[9];
	assign m[10] = ((~( en[10] & en[9] & en[8] )) & s[2]) ^ b[10];
	assign m[11] = ((~( en[11] & en[10] & en[9] )) & s[0]) ^ b[11];
	assign m[12] = ((~( en[12] & en[11] & en[10] )) & s[1]) ^ b[12];
	assign m[13] = ((~( en[13] & en[12] & en[11] )) & s[2]) ^ b[13];
	assign m[14] = ((~( en[14] & en[13] & en[12] )) & s[0]) ^ b[14];
	assign m[15] = ((~( en[15] & en[14] & en[13] )) & s[1]) ^ b[15];
	assign m[16] = ((~( en[16] & en[15] & en[14] )) & s[2]) ^ b[16];
	assign m[17] = ((~( en[17] & en[16] & en[15] )) & s[0]) ^ b[17];
	assign m[18] = ((~( en[18] & en[17] & en[16] )) & s[1]) ^ b[18];
	assign m[19] = ((~( en[19] & en[18] & en[17] )) & s[2]) ^ b[19];
	assign m[20] = ((~( en[20] & en[19] & en[18] )) & s[0]) ^ b[20];
	assign m[21] = ((~( en[21] & en[20] & en[19] )) & s[1]) ^ b[21];
	assign m[22] = ((~( en[22] & en[21] & en[20] )) & s[2]) ^ b[22];
	assign m[23] = ((~( en[23] & en[22] & en[21] )) & s[0]) ^ b[23];
	assign m[24] = ((~( en[24] & en[23] & en[22] )) & s[1]) ^ b[24];
	assign m[25] = ((~( en[25] & en[24] & en[23] )) & s[2]) ^ b[25];
	assign m[26] = ((~( en[26] & en[25] & en[24] )) & s[0]) ^ b[26];
	assign m[27] = ((~( en[27] & en[26] & en[25] )) & s[1]) ^ b[27];
	assign m[28] = ((~( en[28] & en[27] & en[26] )) & s[2]) ^ b[28];
	assign m[29] = ((~( en[29] & en[28] & en[27] )) & s[0]) ^ b[29];
	assign m[30] = ((~( en[30] & en[29] & en[28] )) & s[1]) ^ b[30];
	assign m[31] = ((~( en[31] & en[30] & en[29] )) & s[2]) ^ b[31];

endmodule